`include "uvm_macros.svh"
`include "jtag_pkg.sv"
`include "jtag_if.sv"

//------------------------------------------------------------------------------
// Module: system_shell
//   This is the DUT.
//------------------------------------------------------------------------------

module system_shell( jtag_if.slave_mp jtag_if );
   import jtag_pkg::*;
  
   
endmodule: system_shell

